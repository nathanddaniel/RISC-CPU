
module DataPath(

  //control signals for outputting data to the bus
  input PCout, Zhighout, Zlowout, MDRout, BAout, Rin, Rout,
  input HIout, LOout, Yout, InPortout, Cout, OutPortin,

  //control signals for writing to registers
  input MARin, PCin, MDRin, IRin, Yin, CONin,
  input IncPC, Read, Write,

  //register selection and instruction decoding
	input Gra, Grb, Grc, 				 
  input [4:0] opcode,
  input HIin, LOin, ZHighIn, ZLowIn,

  //global signals
  input clock, clear,

  //address for memory access
  input [8:0] Address,

  //data from memory
  input [31:0] Mdatain,

  //external input
	input wire [31:0] InPortData,
	 
  //outputs from the general registers and OutPort
	output R0out, R1out, R2out, R3out, R4out, R5out, R6out, R7out,
  output R8out, R9out, R10out, R11out, R12out, R13out, R14out, R15out,

  //output to external port
	output wire [31:0] OutPortData

);

//ALU output to the Z regiser
wire [63:0] BusMuxInZ;

//bus inputs from the general regisetrs as well as the special-purpose registers
wire [31:0] BusMuxInR0, BusMuxInR1, BusMuxInR2, BusMuxInR3;
wire [31:0] BusMuxInR4, BusMuxInR5, BusMuxInR6, BusMuxInR7;
wire [31:0] BusMuxInR8, BusMuxInR9, BusMuxInR10, BusMuxInR11;
wire [31:0] BusMuxInR12, BusMuxInR13, BusMuxInR14, BusMuxInR15;
wire [31:0] BusMuxInHI, BusMuxInLO, BusMuxInY;
wire [31:0] BusMuxInZhigh, BusMuxInZlow;
wire [31:0] BusMuxInPC, BusMuxInMDR, BusMuxIn_InPort, BusMuxInCsignextended;

//final bus output
wire [31:0] BusMuxOut;

//memory and bus signals  
wire [8:0]  mem_address;
wire [31:0] mem_data_out;
wire [31:0] mem_data_in;

//signals generated by select and encode logic
wire [15:0] RinSignals, RoutSignals;

//direct output of the MDR
wire [31:0] MDR_data_out;

//IR and instruction decoding 
wire [31:0] IR_out;
wire [4:0] Opcode;
wire [3:0] Ra, Rb, Rc;
wire [18:0] C;
wire [3:0] C2;
wire CON_out;
  

//instantiating the register R0
r0 r0_inst (
	.clear(clear), .clock(clock), .enable(R0in),
	.BAout(BAout), .BusMuxOut(BusMuxOut), .BusMuxIn(BusMuxInR0)
);
	
//the rest of the register instantiations
register r1 (clear, clock, R1in,  BusMuxOut, BusMuxInR1);
register r2 (clear, clock, R2in,  BusMuxOut, BusMuxInR2);
register r3 (clear, clock, R3in,  BusMuxOut, BusMuxInR3);
register r4 (clear, clock, R4in,  BusMuxOut, BusMuxInR4);
register r5 (clear, clock, R5in,  BusMuxOut, BusMuxInR5);
register r6 (clear, clock, R6in,  BusMuxOut, BusMuxInR6);
register r7 (clear, clock, R7in,  BusMuxOut, BusMuxInR7);
register r8 (clear, clock, R8in,  BusMuxOut, BusMuxInR8);
register r9 (clear, clock, R9in,  BusMuxOut, BusMuxInR9);
register r10 (clear, clock, R10in, BusMuxOut, BusMuxInR10);
register r11 (clear, clock, R11in, BusMuxOut, BusMuxInR11);
register r12 (clear, clock, R12in, BusMuxOut, BusMuxInR12);
register r13 (clear, clock, R13in, BusMuxOut, BusMuxInR13);
register r14 (clear, clock, R14in, BusMuxOut, BusMuxInR14);
register r15 (clear, clock, R15in, BusMuxOut, BusMuxInR15);

//special-purpose registers
register HI (clear, clock, HIin,  BusMuxOut, BusMuxInHI);
register LO (clear, clock, LOin,  BusMuxOut, BusMuxInLO);
register Y (clear, clock, Yin,   BusMuxOut, BusMuxInY);
register Zhigh (clear, clock, ZHighIn, BusMuxInZ[63:32], BusMuxInZhigh);
register Zlow (clear, clock, ZLowIn,  BusMuxInZ[31:0],  BusMuxInZlow);
  
//instantiating the CONFF logic
CON_FF con_ff (
  .Clock(clock), .Clear(clear), .CONin(CONin), 
  .BusMuxOut(BusMuxOut), .C2(C2), .CON(CON_out)           
);

//instantiating the program counter logic
ProgramCounter PC_inst (
	.clock(clock), .clear(clear), .enable(PCin), .IncPC(IncPC), .CON(CON_out),                              
	.inputPC(BusMuxOut), .C_sign_extended(BusMuxInCsignextended), .newPC(BusMuxInPC)                      
);
  
//assigning register enable signals (both RXin and RYout, where X and Y represent integers from 0-15)
assign {R15in, R14in, R13in, R12in, R11in, R10in, R9in, R8in, 
        R7in, R6in, R5in, R4in, R3in, R2in, R1in, R0in} = RinSignals;

assign {R15out, R14out, R13out, R12out, R11out, R10out, R9out, R8out, 
        R7out, R6out, R5out, R4out, R3out, R2out, R1out, R0out} = RoutSignals;  
  
//instantiating the Memory Address register
MAR mar_inst (
  .BusMuxOut(BusMuxOut), .MARin(MARin), .Clock(clock), 
  .Clear(clear), .Address(mem_address) //connecting to the RAM
);
  
//instantiating the RAM 
RAM ram_inst (
  .Read(Read), .Write(Write), .Clock(clock), 
  .Mdatain(BusMuxOut), .Address(mem_address), 
  .data_output(mem_data_out) //output to MDR
);
  
//instantiating the Memory Data Register
mdr mdr_inst (
  .Clear(clear), .Clock(clock), .MDRin(MDRin), 
  .Read(Read), .BusMuxOut(BusMuxOut), 
  .Mdatain(mem_data_out), //data from RAM
  .BusMuxIn(BusMuxInMDR), //output to CPU Bus
	.MDR_data_out(MDR_data_out)
);
  
  
//Bus Mux instantiation
Bus bus (
  .BusMuxInR0(BusMuxInR0), .BusMuxInR1(BusMuxInR1), .BusMuxInR2(BusMuxInR2), .BusMuxInR3(BusMuxInR3),
  .BusMuxInR4(BusMuxInR4), .BusMuxInR5(BusMuxInR5), .BusMuxInR6(BusMuxInR6), .BusMuxInR7(BusMuxInR7),
  .BusMuxInR8(BusMuxInR8), .BusMuxInR9(BusMuxInR9), .BusMuxInR10(BusMuxInR10), .BusMuxInR11(BusMuxInR11),
  .BusMuxInR12(BusMuxInR12), .BusMuxInR13(BusMuxInR13), .BusMuxInR14(BusMuxInR14), .BusMuxInR15(BusMuxInR15),
  .BusMuxInHI(BusMuxInHI), .BusMuxInLO(BusMuxInLO), .BusMuxInY(BusMuxInY), .BusMuxInZhigh(BusMuxInZhigh),
  .BusMuxInZlow(BusMuxInZlow), .BusMuxInPC(BusMuxInPC), .BusMuxInMDR(BusMuxInMDR),
  .BusMuxIn_InPort(BusMuxIn_InPort), .BusMuxInCsignextended(BusMuxInCsignextended),

  .PCout(PCout), .Zhighout(Zhighout), .Zlowout(Zlowout), .MDRout(MDRout),
  .R0out(R0out), .R1out(R1out), .R2out(R2out), .R3out(R3out), .R4out(R4out), .R5out(R5out), 
  .R6out(R6out), .R7out(R7out), .R8out(R8out), .R9out(R9out), .R10out(R10out), .R11out(R11out), 
  .R12out(R12out), .R13out(R13out), .R14out(R14out), .R15out(R15out), 
  .HIout(HIout), .LOout(LOout), .Yout(Yout), .InPortout(InPortout), .Cout(Cout), .BAout(BAout),

  .BusMuxOut(BusMuxOut)
);

//instantiating the select and encode logic 
select_and_encode selectLogic (
  .Gra(Gra), .Grb(Grb),	.Grc(Grc),
  .Rin(Rin), .Rout(Rout), .BAout(BAout),
  .Ra(Ra), .Rb(Rb), .Rc(Rc), .C(C),       						 
  .RinSignals(RinSignals), .RoutSignals(RoutSignals),    
  .C_sign_extended(BusMuxInCsignextended) 
);
  
//ALU instantiation
ALU main_alu (
	.clear (clear), .clock (clock), .opcode(opcode),
	.A (BusMuxInY), //operand A recieves value from reg Y   
	.B (BusMuxOut), //operand B recieves value from bus  
	.Z (BusMuxInZ) //Result is stored in reg Z
);
  
//IR instantiation
IR ir_inst (
	.Clock(clock), .Clear(clear), .IRin(IRin),
	.BusMuxOut(BusMuxOut), //getting the instruction from bus
	.IR(IR_out), //storing the instruction
	.Opcode(Opcode), //extracting the opcode fieeld
	.Ra(Ra), .Rb(Rb), .Rc(Rc), //extracting the register fields
	.C(C), //extracting the constant field
	.C2(C2), //extracting the branch condition field 
	.Jaddr(Jaddr) //extracting the jump address
);
	
//InPort instantiation
InPort inport_inst (
	.clock(clock), .clear(clear),
	.InPortData(InPortData), //this is the external input signal
	.BusMuxIn_InPort(BusMuxIn_InPort) //connecting to the CPU bus
);

//OutPort instantiation
OutPort outport_inst (
	.clock(clock), .clear(clear),
	.OutPortin(OutPortin), //enable for OutPort
	.BusMuxOut(BusMuxOut), //data from the Bus
	.OutPortData(OutPortData) //connecting to the external output
);

endmodule